module funcs

pub fn banner(){
	println("
╔════════╦══════════════════════════════════╗
║ Menu # ║ Password Manager by WhosGotFrost ║
╠════════╬══════════════════════════════════╣
║ 1.     ║ Add Password                     ║
║ 2.     ║ Your Saved Passwords             ║
║ 3.     ║ Clears Password txt file         ║
║ exit   ║ will exit the tool               ║
╚════════╩══════════════════════════════════╝
	")
}
